module getLCDdata(score, data_bit, write_enable);
	reg char_count;
	output[7:0] data_bit;
	output write_enable;
	
	
	
endmodule;